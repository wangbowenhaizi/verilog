module timer();

endmodule
`timescale 1ns/1ns
module fer_tb();
output clk,en,count_en,count_clr;
wire clk,en,count_en,count_clr;

endmodule